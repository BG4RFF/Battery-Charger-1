plot the result

.control

load rawspice.raw


*User defined vector and plot commands: 

plot zener

.endc 
.end 

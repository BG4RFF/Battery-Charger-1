plot the result

.control

load rawspice.raw


*User defined vector and plot commands: 

plot i(v2) i(vp2) i(vp3) panelm isolate

.endc 
.end 

plot the result

.control

load rawspice.raw


*User defined vector and plot commands: 

plot i(vbattery) linear

.endc 
.end 
